   // PMEM
   input  [1-1:0]    pmem_rst_btn,
   input  [10-1:0]   pmem_pixel_x,
   input  [10-1:0]   pmem_pixel_y,
   output [12-1:0]   pmem_rgb,
