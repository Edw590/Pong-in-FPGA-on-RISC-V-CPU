   // PMEM
   input  [32-1:0]   pmem_sw_input,
   input  [10-1:0]   pmem_pixel_x,
   input  [10-1:0]   pmem_pixel_y,
   output [12-1:0]   pmem_rgb,
