   // IM
   input  [32-1:0]   im_sw_input,
   input  [10-1:0]   im_pixel_x,
   input  [10-1:0]   im_pixel_y,
   input  [8-1:0]    im_ctrl1_data,
   input  [8-1:0]    im_ctrl2_data,
   output [12-1:0]   im_rgb,
