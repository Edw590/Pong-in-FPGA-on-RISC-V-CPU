   // IM
   input  [32-1:0]   im_sw_input,
   input  [10-1:0]   im_pixel_x,
   input  [10-1:0]   im_pixel_y,
   output [12-1:0]   im_rgb,
